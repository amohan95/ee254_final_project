`define X_MAX 640
`define Y_MAX 480