`include "constants.vh"

module vga_controller(input wire clk, reset,
                      input wire [9:0] CounterX, CounterY,
                      output reg [2:0] r, g,
                      output reg [1:0] b);
  
endmodule