module game_controller(input wire clk, reset);
  `include "constants.vh"
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      
    end
    else begin
      
    end
  end
endmodule