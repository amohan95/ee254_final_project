module vga_controller(clk, reset, vga_h_sync, vga_v_sync, inDisplayArea, CounterX, CounterY);